//
// 存放所有 ASCII 字符的字码
// 该ROM自动综合成Block RAM
// 每个字符为8*16个像素，8列16行
// 机制：每次读取时需要输入一个 7bit ASCII 值和一个 4bit 行号，共同组成12bit地址
// ASCII值表示想要读取的字符的ASCII码
// 4bit行号的取值范围是0~15，指定了想要读取该字符的哪一行像素。
// 输出8bit，即该字符这一行的8个像素。0代表黑色，1代表白色（黑底白字）
// 因此该模块只是一个普通的8bit数据总线，12bit地址总线的ROM而已

module char8x16_rom(
    input  logic clk,
    input  logic [11:0] addr,
    output logic [ 7:0] data
);

wire [0:2047] [7:0] rom_cell = {
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h10,
    8'h00,
    8'h10,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h2c,
    8'h24,
    8'h24,
    8'h24,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h68,
    8'h24,
    8'hfe,
    8'h24,
    8'h24,
    8'h24,
    8'h7e,
    8'h24,
    8'h24,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h10,
    8'h7c,
    8'h16,
    8'h12,
    8'h16,
    8'h38,
    8'h68,
    8'h48,
    8'h48,
    8'h3e,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h86,
    8'h4b,
    8'h69,
    8'h2e,
    8'h10,
    8'h08,
    8'h68,
    8'h94,
    8'h92,
    8'h63,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h26,
    8'h26,
    8'h1c,
    8'h4e,
    8'h52,
    8'h73,
    8'h62,
    8'hfe,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h10,
    8'h18,
    8'h08,
    8'h0c,
    8'h0c,
    8'h0c,
    8'h0c,
    8'h08,
    8'h08,
    8'h18,
    8'h30,
    8'h20,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h08,
    8'h10,
    8'h10,
    8'h30,
    8'h20,
    8'h20,
    8'h20,
    8'h30,
    8'h10,
    8'h18,
    8'h08,
    8'h04,
    8'h00,
    8'h00,
    8'h00,
    8'h10,
    8'h50,
    8'h2c,
    8'h38,
    8'h56,
    8'h10,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'hfe,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h10,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h40,
    8'h60,
    8'h20,
    8'h30,
    8'h10,
    8'h10,
    8'h08,
    8'h08,
    8'h04,
    8'h04,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h66,
    8'h42,
    8'he2,
    8'hda,
    8'hce,
    8'h42,
    8'h66,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h1e,
    8'h12,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h62,
    8'h60,
    8'h60,
    8'h20,
    8'h10,
    8'h08,
    8'h04,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h60,
    8'h60,
    8'h20,
    8'h3c,
    8'h40,
    8'h40,
    8'h60,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h30,
    8'h38,
    8'h28,
    8'h24,
    8'h26,
    8'h22,
    8'hff,
    8'h20,
    8'h20,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h40,
    8'h40,
    8'h60,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h0c,
    8'h06,
    8'h12,
    8'h6e,
    8'h42,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h40,
    8'h60,
    8'h20,
    8'h30,
    8'h10,
    8'h18,
    8'h08,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'h6c,
    8'h38,
    8'h66,
    8'h42,
    8'h42,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h66,
    8'h42,
    8'h42,
    8'h66,
    8'h58,
    8'h40,
    8'h20,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h10,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h18,
    8'h0c,
    8'h06,
    8'h08,
    8'h30,
    8'h60,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h00,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h18,
    8'h20,
    8'h60,
    8'h30,
    8'h08,
    8'h04,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h38,
    8'h60,
    8'h60,
    8'h60,
    8'h18,
    8'h08,
    8'h00,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h38,
    8'h44,
    8'h82,
    8'h82,
    8'hbb,
    8'had,
    8'ha5,
    8'ha5,
    8'hf5,
    8'h29,
    8'h03,
    8'h02,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h38,
    8'h2c,
    8'h24,
    8'h64,
    8'h46,
    8'h7e,
    8'hc2,
    8'h83,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'h62,
    8'h3e,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h04,
    8'h02,
    8'h02,
    8'h02,
    8'h02,
    8'h02,
    8'h06,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'hc2,
    8'hc2,
    8'hc2,
    8'h42,
    8'h62,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h06,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h06,
    8'h02,
    8'h02,
    8'h73,
    8'h42,
    8'h42,
    8'h46,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h7e,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h22,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h22,
    8'h12,
    8'h0a,
    8'h0e,
    8'h1a,
    8'h32,
    8'h22,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h66,
    8'he6,
    8'hfa,
    8'hda,
    8'hda,
    8'h83,
    8'h83,
    8'h83,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h46,
    8'h4e,
    8'h4a,
    8'h5a,
    8'h52,
    8'h72,
    8'h62,
    8'h62,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'hc2,
    8'hc3,
    8'hc3,
    8'hc3,
    8'hc2,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'h42,
    8'h62,
    8'h1e,
    8'h02,
    8'h02,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'hc2,
    8'hc3,
    8'hc3,
    8'hc3,
    8'hc2,
    8'h46,
    8'h3c,
    8'h18,
    8'hf0,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h66,
    8'h46,
    8'h66,
    8'h3e,
    8'h36,
    8'h26,
    8'h66,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h06,
    8'h02,
    8'h06,
    8'h38,
    8'h60,
    8'h40,
    8'h40,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hfe,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'hc2,
    8'h42,
    8'h46,
    8'h64,
    8'h24,
    8'h2c,
    8'h38,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h83,
    8'h82,
    8'h92,
    8'hda,
    8'hda,
    8'h6e,
    8'h66,
    8'h66,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h66,
    8'h2c,
    8'h18,
    8'h18,
    8'h38,
    8'h24,
    8'h66,
    8'hc3,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h42,
    8'h66,
    8'h2c,
    8'h38,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h40,
    8'h20,
    8'h30,
    8'h18,
    8'h08,
    8'h04,
    8'h06,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h38,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h38,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h04,
    8'h04,
    8'h08,
    8'h08,
    8'h10,
    8'h10,
    8'h30,
    8'h20,
    8'h60,
    8'h40,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h38,
    8'h24,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hff,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h60,
    8'h40,
    8'h7c,
    8'h42,
    8'h62,
    8'h5e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h02,
    8'h02,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h04,
    8'h06,
    8'h02,
    8'h06,
    8'h04,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h40,
    8'h40,
    8'h40,
    8'h7c,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'h7e,
    8'h02,
    8'h06,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hf0,
    8'h18,
    8'h08,
    8'h08,
    8'h7e,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hfc,
    8'h66,
    8'h42,
    8'h66,
    8'h1a,
    8'h02,
    8'h7c,
    8'hc2,
    8'h42,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h02,
    8'h02,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h1e,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h30,
    8'h00,
    8'h3e,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h30,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h06,
    8'h06,
    8'h06,
    8'h46,
    8'h36,
    8'h1e,
    8'h0e,
    8'h16,
    8'h26,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h1e,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h6e,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'hc2,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h02,
    8'h02,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h40,
    8'h40,
    8'h40,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h76,
    8'h4e,
    8'hc6,
    8'h06,
    8'h06,
    8'h06,
    8'h06,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h04,
    8'h04,
    8'h3c,
    8'h60,
    8'h40,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h08,
    8'h08,
    8'h7f,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h78,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h42,
    8'h66,
    8'h24,
    8'h2c,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h83,
    8'hda,
    8'h5a,
    8'h7a,
    8'h66,
    8'h66,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h64,
    8'h38,
    8'h18,
    8'h38,
    8'h64,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h42,
    8'h66,
    8'h24,
    8'h2c,
    8'h38,
    8'h18,
    8'h18,
    8'h0c,
    8'h07,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h60,
    8'h30,
    8'h18,
    8'h08,
    8'h04,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h70,
    8'h18,
    8'h08,
    8'h08,
    8'h08,
    8'h0c,
    8'h0e,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h18,
    8'h70,
    8'h00,
    8'h00,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h18,
    8'h10,
    8'h10,
    8'h10,
    8'h30,
    8'h70,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h18,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h8e,
    8'hd2,
    8'h60,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00
};

always @ (posedge clk)
    if(addr[11])
        data <= 8'h0;
    else
        data <= rom_cell[addr[10:0]];

endmodule
